----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:31:50 05/09/2020 
-- Design Name: 
-- Module Name:    T_FF - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity T_FF is
    Port ( CLK : in  STD_LOGIC;
           T : in  STD_LOGIC;
           Q : out  STD_LOGIC;
           Qn : out  STD_LOGIC);
end T_FF;

architecture Behavioral of T_FF is

signal temp, tempn:STD_LOGIC:='0';

begin
	process(CLK, T)
	begin
		if rising_edge(CLK) then
			if T = '0' then
				temp <= temp;
				tempn <= tempn;
			else
				temp <= not temp;
				tempn <= not tempn;
			end if;
		end if;
	end process;
Q<=temp; Qn<=tempn;
end Behavioral;

